module board (
  input logic CLK, RST
);

endmodule // board
